000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111111111111111111111111111111000111111111111111111111111110001111111111111111111111111100111111111111111111111111111111001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000001111111111111111111111111111111000111111111111111111111111110001111111111111111111111111100111111111111111111111111111111001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000001111111111111111111111111111111000111111111111111111111111110001111111111111111111111111100111111111111111111111111111111001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000001111111111111111111111111111111000111111111111111111111111110001111111111111111111111111100111111111111111111111111111111001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000000000111100000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000000001111000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000000011110000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000000111100000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000001111000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000011110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000000111100000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000001111000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000011110000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000000111100000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000000000000000000000001111000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111111111111111111111111110001111000000000000000000111100000000000000011111000000000000000000000000000000011110000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111111111111111111111111110001111000000000000000000111100000000000000011111000000000000000000000000000000111100000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111111111111111111111111110001111000000000000000000111100000000000000011111000000000000000000000000000001111000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000011111000000000001111000000000000000000111100000000000000011111000000000000000000000000000011110000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000001111000000000001111111111111111111111111100000000000000011111000000000000000000000000000111100000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000000000000111100000000000111100000000001111111111111111111111111100000000000000011111000000000000000000000000001111000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000001111111111111000111100000000000111100000000001111111111111111111111111100000000000000011111000000000000000000000000011110000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000001111111111111000111100000000000011110000000001111000000000000000000111100000000000000011111000000000000000000000000111100000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000001111111111111000111100000000000011110000000001111000000000000000000111100000000000000011111000000000000000000000001111000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000001111111111111000111100000000000001111000000001111000000000000000000111100000000000000011111000000000000000000000011110000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000001111000000001111000000000000000000111100000000000000011111000000000000000000000111100000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000111100000001111000000000000000000111100000000000000011111000000000000000000001111000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000111100000001111000000000000000000111100000000000000011111000000000000000000011110000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000011110000001111000000000000000000111100000000000000011111000000000000000000111100000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000011110000001111000000000000000000111100000000000000011111000000000000000001111000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000001111000001111000000000000000000111100000000000000011111000000000000000011110000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000001111000001111000000000000000000111100000000000000011111000000000000000111100000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000111100000000000000000111100001111000000000000000000111100000000000000011111000000000000001111100000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111111111111111111111111111111000111100000000000000000111100001111000000000000000000111100000000000000011111000000000000001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000000111111111111111111111111111110000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000000011111111111111111111111111100000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000000001111111111111111111111111000000111100000000000000000011110001111000000000000000000111100000000000000011111000000000000001111111111111111111111111111111110000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111111111111111111111000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111111111111111111111100000000001111111111111111111111111100000000000000000000000000000000000000000010000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111111111111111111111110000000001111111111111111111111111100000000000000000000000000000000000011000010000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111111111111111111111111000000001111111111111111111111111100000000000000000000000000000000010001000110000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000111100000001111000000000000000000111100000000000000000000000000000000001001001000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000011110000001111000000000000000000111100000000000000000000000000000000000101010000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000001111000001111000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000111100001111000000000000000000111100000000000000000000000000000000000011001111110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000011111001111000000000000000000111100000000000000000000000000000000000011001000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000000000000000001100001000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000000000000000011000000100000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000000000000000110000000100000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000000000000001100000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000000000000001100000000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000000000001111111110000000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111111111111111111111111100000000000000000000000000111111111111100000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111111111111111111111111100000000000000000000000001111111111111110000000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111111111111111111111111100000000000000000000000111111111111111111100000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000001111111111111111111110000000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000000111111111111111111111111100000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000001111111111111111111111111110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000001111111111111111111111111110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000001111001111000000000000000000111100000000000000000001111111111111111111111111110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000011110001111000000000000000000111100000000000000000001111111111111111111111111110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000000111100001111000000000000000000111100000000000000000001111111111111111111111111110000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000001111000001111000000000000000000111100000000000000000000111111111111111111111111100000000000000000000000000000000
000000000000000000000000000000001111000000000000000000000001111000000000000000111100000000000000000011110000001111000000000000000000111100000000000000000000001111111111111111111110000000000000000000000000000000000
000000000000000000000000000000001111111111111111111111111111111000000000000000111111111111111111111111000000001111000000000000000000111100000000000000000000000111111111111111111100000000000000000000000000000000000
000000000000000000000000000000000111111111111111111111111111110000000000000000111111111111111111111110000000001111000000000000000000111100000000000000000000000001111111111111110000000000000000000000000000000000000
000000000000000000000000000000000011111111111111111111111111100000000000000000111111111111111111111100000000001111000000000000000000111100000000000000000000000000111111111111100000000000000000000000000000000000000
000000000000000000000000000000000001111111111111111111111111000000000000000000111111111111111111111000000000001111000000000000000000111100000000000000000000000000001111111110000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000


