00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111111111111111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111111111111111111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000011111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000001111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000111111000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111100000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000011111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000001111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111111111111000000000000000000000000000111111111111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111000000000000000000000111111000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111111111110000000000000000001111111110000000001111111110000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111000000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111100000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111110000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000011111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000001111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000111111111000000000000000000000111111000000000000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111000000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111100000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111110000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000010001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000011111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000001111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111000000000000000000111111111000000000000000000000111111000000000000000000000000000111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111000000000000000000000111111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111100000000000000000000111111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111110000000000000000000111111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000111111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000011111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000001111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000111111111111111111111111111111111000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000111111111000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000111111111000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000111111111000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000111111111000000000000000001111111110000000000000000001111111110000000001111111110000000000000000001111111110000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
11111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111110000000001111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
