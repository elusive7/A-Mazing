0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111111111111100000000000000000000000000000000000000000000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111100000000011111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111111111111111111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111111111111111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000001111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000111111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000011111100000000000000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111100000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111110000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000001111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000000111111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111111111111100000000000000000000000000011111111111111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111100000000000000000000011111100000000000000000000000000000000000000000000011111111100000000000000000011111111111111111111111111111111111000000000000000000111111111000000000111111111000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111100000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111110000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111000000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000001111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000000111111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000011111111100000000000000000000011111100000000000000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111100000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111110000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111000000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000001000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111100000000000000000001111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000111111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
0000000011111111100000000011111111100000000000000000011111111100000000000000000011111111100000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111100000000000000000011111111100000000000000000000011111100000000000000000000000000011111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111100000000000000
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111100000000000000000000011111111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111110000000000000000000011111111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111000000000000000000011111111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000011111111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000001111111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000111111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000011111111111111111111111111111111111111111111100000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000011111111111111111111111111111111100000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
1111111111111111100000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000011111111100000000000000000011111111111111111111111
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
0000000000000000000000000011111111100000000000000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000011111111100000000000000000000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000011111111100000000000000000111111111000000000000000000111111111000000000111111111000000000000000000111111111000000000000000011111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000011111111100000000000000000000000000000000000000000
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111
1111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111000000000111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111

