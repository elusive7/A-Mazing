00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000001'b1,0001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,000000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,00000000000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000001'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000

