1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1'b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,
1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1'b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b1,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,1’b0,

